// Generate by chisel-memory-lower
// Target: arm
// Config(name='mem_1rw', depth='48', width='64', ports='rw', mask_gran=None)
module mem_1rw (
  input [5:0] RW0_addr,
  input RW0_en,
  input RW0_clk,
  input RW0_wmode,
  input [63:0] RW0_wdata,
  output [63:0] RW0_rdata
);

endmodule
