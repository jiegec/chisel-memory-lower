// Generate by chisel-memory-lower
// Target: arm
// Config(name='mem_1r1w', depth='32', width='64', ports='write,read', mask_gran=None)
module mem_1r1w (
  input [4:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [63:0] R0_data,
  input [4:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [63:0] W0_data
);

endmodule
